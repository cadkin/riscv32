`timescale 1ns/1ps

module fcsr();
	// foobar
endmodule;
